----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:17:08 04/08/2019 
-- Design Name: 
-- Module Name:    ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_unsigned.ALL ;
use IEEE.std_logic_arith.ALL ;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ROM is
	port (
			Address : in std_logic_vector ( 9 downto 0 ) ;
			Data_out : out std_logic_vector ( 15 downto 0 ) );
end ROM;

architecture Behavioral of ROM is

type ram is array ( 0 to(2**12) ) of std_logic_vector ( 15 downto 0 ) ;
constant in_reg : ram := 
("0000000000000001",
"0100000000010000",
"0000000000000110",
"0010000000000000",
"0000110110110001",
"0000001001001001",
"0100110110011111",
"0100110110010100",
"1000110001000000",
"0000110110110001",
"0100110110001001",
"1000110001000000",
"0000100100100001",
"1100000101100011",
"0000110110110001",
"0100110110001001",
"0111110010000000",
"0000001001001001",
"0100001001000001",
"1001010001000001",
"1011000000001101",
"0000010010010001",
"1000110010000000",
"0000110110110001",
"0100110110001000",
"0111110010000000",
"0000001001001001",
"0000010000010111",
"1001010001000001",
"1011000000100000",
"0100100100010100",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000000100101",
"0100100100011001",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000000101010",
"0100100100001111",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000000101111",
"0100100100011110",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000000110100",
"0100100100011001",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000000111001",
"0100100100011001",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000000111110",
"0100100100010100",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000001000011",
"0100100100001010",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000001001000",
"0100100100001111",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000001001101",
"0100100100010100",
"1011000000001101",
"0000010000010111",
"1001010001000001",
"1011000000001101",
"0000110110110001",
"0100110110001110",
"1000110100000000",
"1100000101100011",
"0000110110110001",
"0100110110001001",
"0111110010000000",
"0000001001001001",
"0100001001000001",
"1001010001000001",
"1011000001010011",
"1011000000001100",
"1110000000000000",
"0000110110110001",
"1000110000000000",
"0100110110000001",
"1000110001000000",
"0100110110000001",
"1000110010000000",
"0100110110000001",
"1000110011000000",
"0100110110000001",
"1000110100000000",
"0100110110000001",
"1000110101000000",
"0000001001001001",
"0000110110110001",
"0100110110001101",
"0000010010010001",
"0111110010000000",
"0000010001001011",
"0010001000000000",
"0000011011011001",
"0100011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0110011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000100100100001",
"0000101101101001",
"0100101101000001",
"1001011100000010",
"0000011101011001",
"1011000001111111",
"0000010010010001",
"0100010010000001",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010001001011",
"0010001000000000",
"0000011011011001",
"0100011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0110011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000100100100001",
"0000101101101001",
"0100101101000001",
"1001011100000010",
"0000011101011001",
"1011000010011101",
"0000010010010001",
"0100010010011111",
"0100010010011111",
"0100010010011111",
"0100010010011111",
"0100010010011111",
"0100010010011111",
"0100010010011111",
"0100010010011111",
"0100010010000111",
"0000001010001010",
"0010001000000000",
"0000011011011001",
"0100011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0110011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000100100100001",
"0000101101101001",
"0100101101000001",
"1001011100000010",
"0000011101011001",
"1011000010111011",
"0000110110110001",
"0111110000000000",
"0100110110000001",
"0111110001000000",
"0100110110000001",
"0111110010000000",
"0100110110000001",
"0111110011000000",
"0100110110000001",
"0111110100000000",
"0100110110000001",
"0111110101000000",
"0011111000000000",
"1110000000000000",
"0000110110110001",
"1000110000000000",
"0100110110000001",
"1000110001000000",
"0100110110000001",
"1000110010000000",
"0100110110000001",
"1000110011000000",
"0100110110000001",
"1000110100000000",
"0100110110000001",
"1000110101000000",
"0000001001001001",
"0100001001000001",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000110110110001",
"0100110110001100",
"0000010010010001",
"0111110010000000",
"0000010001001011",
"0010001000000000",
"0000011011011001",
"0100011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0110011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000100100100001",
"0000101101101001",
"0100101101000001",
"1001011100000010",
"0000011101011001",
"1011000011111000",
"0000010010010001",
"0100010010000001",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010001001011",
"0010001000000000",
"0000011011011001",
"0100011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0110011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000100100100001",
"0000101101101001",
"0100101101000001",
"1001011100000010",
"0000011101011001",
"1011000100010110",
"0000010010010001",
"0100010010010111",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000010000010110",
"0000011011011001",
"0100011011011111",
"0000011010010011",
"0000001010001010",
"0010001000000000",
"0000011011011001",
"0100011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0110011011011111",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000011000011110",
"0000100100100001",
"0000101101101001",
"0100101101000001",
"1001011100000010",
"0000011101011001",
"1011000100110100",
"0000110110110001",
"0111110000000000",
"0100110110000001",
"0111110001000000",
"0100110110000001",
"0111110010000000",
"0100110110000001",
"0111110011000000",
"0100110110000001",
"0111110100000000",
"0100110110000001",
"0111110101000000",
"0011111000000000",
"1110000000000000",
"0000110110110001",
"1000110000000000",
"0000110110110001",
"0100110110000111",
"1000110111000000",
"0000000000000001",
"0100000000011110",
"0100000000011010",
"0000110110110001",
"0100110110001101",
"1000110000000000",
"1100000001011100",
"0000000000000001",
"0100000000001100",
"0000110110110001",
"0100110110001101",
"1000110000000000",
"1100000001011100",
"0000000000000001",
"0100000000000001",
"0000110110110001",
"0100110110001101",
"1000110000000000",
"1100000001011100",
"0000110110110001",
"0111110000000000",
"0000110110110001",
"0100110110000111",
"0111110111000000",
"0011111000000000",
"0000110110110001",
"1000110000000000",
"0100110110000001",
"1000110001000000",
"0100110110000001",
"1000110010000000",
"0100110110000001",
"1000110011000000",
"0100110110000001",
"1000110100000000",
"0100110110000001",
"1000110101000000",
"0000110110110001",
"0100110110001001",
"0111110000000000",
"0000001001001001",
"1001001000000001",
"1011001011000111",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0111110000000000",
"0000001001001001",
"1010001000000001",
"1011000110001110",
"0000001001001001",
"0100001001000001",
"1010001000000001",
"1011001000011010",
"0000001001001001",
"0100001001000010",
"1010001000000001",
"1011001001111100",
"0000001001001001",
"0100001001000011",
"1010001000000001",
"1011001010011010",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0000001001001001",
"1000110001000000",
"1011000101101111",
"0000100100100001",
"0100100100001111",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0010100000000000",
"0001000000011000",
"0000101101101001",
"1010011101000110",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0000000000000001",
"1000110000000000",
"1011001000011001",
"0000010010010001",
"0000100100100001",
"0100100100000001",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0000100000100110",
"0010100000000000",
"0001000000011000",
"0000101101101001",
"1001011101010011",
"0000110110110001",
"0100110110011111",
"0100110110010101",
"1000110100000000",
"0000110110110001",
"0100110110011111",
"0100110110010110",
"1000110011000000",
"0000000000000001",
"0100000000000001",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"1000110000000000",
"0000110110110001",
"0100110110011111",
"0100110110010111",
"1000110010000000",
"1011001000011001",
"0100010010000001",
"0000100000100111",
"0010100000000000",
"0001000000011000",
"0000101101101001",
"1001011101010011",
"0000110110110001",
"0100110110011111",
"0100110110010101",
"1000110100000000",
"0000110110110001",
"0100110110011111",
"0100110110010110",
"1000110011000000",
"0000000000000001",
"0100000000000001",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"1000110000000000",
"0000110110110001",
"0100110110011111",
"0100110110010111",
"1000110010000000",
"1011001000011001",
"0100010010000001",
"0000100000100111",
"0010100000000000",
"0001000000011000",
"0000101101101001",
"1001011101010011",
"0000110110110001",
"0100110110011111",
"0100110110010101",
"1000110100000000",
"0000110110110001",
"0100110110011111",
"0100110110010110",
"1000110011000000",
"0000000000000001",
"0100000000000001",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"1000110000000000",
"0000110110110001",
"0100110110011111",
"0100110110010111",
"1000110010000000",
"1011001000011001",
"0100010010000001",
"0000100000100111",
"0010100000000000",
"0001000000011000",
"0000101101101001",
"1001011101010010",
"0000110110110001",
"0100110110011111",
"0100110110010101",
"1000110100000000",
"0000110110110001",
"0100110110011111",
"0100110110010110",
"1000110011000000",
"0000000000000001",
"0100000000000001",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"1000110000000000",
"0000110110110001",
"0100110110011111",
"0100110110010111",
"1000110010000000",
"1011000101101111",
"0000000000000001",
"0100000000001111",
"0000000000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000000001000011",
"0000000000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000000001000011",
"0100000001000000",
"0000010010010001",
"0100010010000100",
"0000100100100001",
"0100100100000001",
"0000110110110001",
"0100110110011111",
"0100110110010101",
"0111110000000000",
"0000110110110001",
"0100110110011111",
"0100110110010110",
"0111110001000000",
"0010000000000000",
"0001000000011000",
"1001001011000110",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0000100100100001",
"1000110100000000",
"1011001001111011",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0000100100100001",
"0100100100000010",
"1000110100000000",
"0000101101101001",
"0100101101001000",
"1010101001000111",
"0000110110110001",
"0100110110011111",
"0100110110011000",
"0000100100100001",
"0100100100000000",
"1000110100000000",
"1011001001101010",
"0000101000101111",
"1010101001000111",
"0000110110110001",
"0100110110011111",
"0100110110011000",
"0000100100100001",
"0100100100000001",
"1000110100000000",
"1011001001101010",
"0000101000101111",
"1010101001000111",
"0000110110110001",
"0100110110011111",
"0100110110011000",
"0000100100100001",
"0100100100000010",
"1000110100000000",
"1011001001101010",
"0000101000101111",
"1010101001000110",
"0000110110110001",
"0100110110011111",
"0100110110011000",
"0000100100100001",
"0100100100000011",
"1000110100000000",
"0000110110110001",
"0100110110011111",
"0100110110010111",
"0111110101000000",
"0000101000000110",
"0000000000000110",
"0000000100000000",
"0100000000000001",
"0000110110110001",
"0100110110011111",
"0100110110011001",
"1000110000000000",
"0000110110110001",
"0100110110001001",
"0000000000000001",
"0100000000000001",
"1000110000000000",
"1011000101101111",
"0000110110110001",
"0100110110011111",
"0100110110010101",
"0111110000000000",
"0000110110110001",
"0100110110011111",
"0100110110010110",
"0111110001000000",
"0010000000000000",
"0001000000011000",
"1001001011000111",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0000100100100001",
"0100100100000011",
"1000110100000000",
"1011001010011001",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0000100100100001",
"0100100100000010",
"1000110100000000",
"0000110110110001",
"0100110110001001",
"0000000000000001",
"0100000000000001",
"1000110000000000",
"1011000101101111",
"0000000000000001",
"0100000000001111",
"0000000000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000000001000011",
"0000000000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000000001000011",
"0100000001000000",
"0000010010010001",
"0100010010000100",
"0000100100100001",
"0100100100000001",
"0000110110110001",
"0100110110011111",
"0100110110010101",
"0111110000000000",
"0000110110110001",
"0100110110011111",
"0100110110010110",
"0111110001000000",
"0010000000000000",
"0001000000011000",
"1001001011000110",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0000100100100001",
"1000110100000000",
"1011001011000110",
"0000110110110001",
"0100110110011111",
"0100110110010100",
"0000100100100001",
"0100100100000010",
"1000110100000000",
"1011000101101111",
"0000110110110001",
"0100110110011111",
"0100110110011001",
"0111110000000000",
"0000110110110001",
"0100110110001000",
"0000001001001001",
"0100001001000001",
"0000010010010001",
"0100010010000001",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010000010",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010000011",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010000101",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010000110",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010000111",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010001001",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010001010",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010001011",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010001110",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000010010010001",
"0100010010000100",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000001000001110",
"0000010010010001",
"0100010010001111",
"1010000010000010",
"1000110001000000",
"1011001100011111",
"0000110110110001",
"0100110110001001",
"0000011011011001",
"1000110011000000",
"1011000101101111",
"0000110110110001",
"0111110000000000",
"0100110110000001",
"0111110001000000",
"0100110110000001",
"0111110010000000",
"0100110110000001",
"0111110011000000",
"0100110110000001",
"0111110100000000",
"0100110110000001",
"0111110101000000",
"0011111000000000",
 others => "1110000000000000"
 );

begin
				Data_out <= in_reg(conv_integer(unsigned(Address))) ;
end Behavioral;

